`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:58:20 11/21/2016 
// Design Name: 
// Module Name:    vga_control_module 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`include "vga_params.v"

module vga_control_module3
(
	input VGA_CLK,
	//input[1:0] switch, //added by me
	input [`P_WIDTH-1:0] X, Y, //11 bits in size
	input valid,
	input [44:0] seq1,
	input [44:0] seq2,
	input [3:0] index10,
	input [3:0] index1,
	output [`D_WIDTH-1:0] VGA_R, VGA_G, VGA_B
);
//wire [3:0] index10, index1;
//assign index10 = 4'd3;
//assign index1 = 4'd4;
//reg arrow;
//assign arrow = 1;
//wire [44:0]seq1,seq2;
//assign seq2=45'b010000100001000010000100001000010000100001000;
//assign seq1=45'b000001010111000000011010111011111000001011000;
//assign seq2=45'b000001010111000000011010111011111000001011000;
/*reg rectangle;
always @ (posedge VGA_CLK)
	if(X > 100 && X < `H_ACT-100 && Y > 100 && Y < `V_ACT-100)
		rectangle <= 1'b0;
	else
		rectangle <= 1'b1;

assign VGA_R = valid && rectangle ? `D_WIDTH'b0000 : `D_WIDTH'b0;
assign VGA_G = valid && rectangle ? `D_WIDTH'b0000 : `D_WIDTH'b0;
assign VGA_B = valid && rectangle ? `D_WIDTH'b1111 : `D_WIDTH'b0;*/
reg [11:0] colouroutput;
always @ (posedge VGA_CLK) begin
	if (~valid)begin
		colouroutput <= 0;
	end
	else begin
		if ((index10==4'd0) && (((X>20&&X<30)&&(Y>90&&Y<140)) || ((X>20&&X<50)&&(Y>90&&Y<100)) || ((X>40&&X<50)&&(Y>90&&Y<140)) || ((X>20&&X<50)&&(Y>130&&Y<140)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index10==4'd1) && (((X>35&&X<45)&&(Y>90&&Y<140))  ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index10==4'd2) && (((X>20&&X<50)&&(Y>90&&Y<100)) || ((X>40&&X<50)&&(Y>90&&Y<120)) || ((X>20&&X<50)&&(Y>110&&Y<120)) || ((X>20&&X<30)&&(Y>110&&Y<140)) || ((X>20&&X<50)&&(Y>130&&Y<140)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index10==4'd3) && (((X>20&&X<50)&&(Y>90&&Y<100)) || ((X>40&&X<50)&&(Y>90&&Y<140)) || ((X>20&&X<50)&&(Y>110&&Y<120)) || ((X>20&&X<50)&&(Y>130&&Y<140)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index10==4'd4) && (((X>20&&X<30)&&(Y>90&&Y<120)) || ((X>20&&X<50)&&(Y>110&&Y<120)) || ((X>40&&X<50)&&(Y>90&&Y<140)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end	
		else if ((index10==4'd5) && (((X>20&&X<50)&&(Y>90&&Y<100)) || ((X>20&&X<30)&&(Y>90&&Y<120)) || ((X>20&&X<50)&&(Y>110&&Y<120)) || ((X>40&&X<50)&&(Y>110&&Y<140)) || ((X>20&&X<50)&&(Y>130&&Y<140)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index10==4'd6) && (((X>20&&X<50)&&(Y>90&&Y<100)) || ((X>20&&X<30)&&(Y>90&&Y<140)) || ((X>20&&X<50)&&(Y>110&&Y<120)) || ((X>20&&X<50)&&(Y>130&&Y<140)) || ((X>40&&X<50)&&(Y>110&&Y<140)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
      else if ((index10==4'd7) && ( ((X>20&&X<50)&&(Y>90&&Y<100))&&((X>40&&X<50)&&(Y>90&&Y<140))  ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index10==4'd8) && (((X>20&&X<30)&&(Y>90&&Y<140)) || ((X>20&&X<50)&&(Y>90&&Y<100)) || ((X>40&&X<50)&&(Y>90&&Y<140)) || ((X>20&&X<50)&&(Y>130&&Y<140)) || ((X>20&&X<50)&&(Y>110&&Y<120)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index10==4'd9) && (((X>20&&X<30)&&(Y>90&&Y<120)) || ((X>20&&X<50)&&(Y>90&&Y<100)) || ((X>40&&X<50)&&(Y>90&&Y<140)) || ((X>20&&X<50)&&(Y>110&&Y<120))  ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		//////////////////%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%/////////////////////
		else if ((index1==4'd0) && (((X>60&&X<70)&&(Y>90&&Y<140)) || ((X>60&&X<90)&&(Y>90&&Y<100)) || ((X>80&&X<90)&&(Y>90&&Y<140)) || ((X>60&&X<90)&&(Y>130&&Y<140)) ))begin
			colouroutput[11:0] <=12'b000011111111;
		end
		else if ((index1==4'd1) && (((X>75&&X<85)&&(Y>90&&Y<140))  ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index1==4'd2) && (((X>60&&X<90)&&(Y>90&&Y<100)) || ((X>80&&X<90)&&(Y>90&&Y<120)) || ((X>60&&X<90)&&(Y>110&&Y<120)) || ((X>60&&X<70)&&(Y>110&&Y<140)) || ((X>60&&X<90)&&(Y>130&&Y<140)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index1==4'd3) && (((X>60&&X<90)&&(Y>90&&Y<100)) || ((X>80&&X<90)&&(Y>90&&Y<140)) || ((X>60&&X<90)&&(Y>110&&Y<120)) || ((X>60&&X<90)&&(Y>130&&Y<140)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index1==4'd4) && (((X>60&&X<70)&&(Y>90&&Y<120)) || ((X>60&&X<90)&&(Y>110&&Y<120)) || ((X>80&&X<90)&&(Y>90&&Y<140)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end	
		else if ((index1==4'd5) && (((X>60&&X<90)&&(Y>90&&Y<100)) || ((X>60&&X<70)&&(Y>90&&Y<120)) || ((X>60&&X<90)&&(Y>110&&Y<120)) || ((X>80&&X<90)&&(Y>110&&Y<140)) || ((X>60&&X<90)&&(Y>130&&Y<140)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index1==4'd6) && (((X>60&&X<90)&&(Y>90&&Y<100)) || ((X>60&&X<70)&&(Y>90&&Y<140)) || ((X>60&&X<90)&&(Y>110&&Y<120)) || ((X>60&&X<90)&&(Y>130&&Y<140)) || ((X>80&&X<90)&&(Y>110&&Y<140)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
      else if ((index1==4'd7) && ( ((X>60&&X<90)&&(Y>90&&Y<100))&&((X>80&&X<90)&&(Y>90&&Y<140))  ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index1==4'd8) && (((X>60&&X<70)&&(Y>90&&Y<140)) || ((X>60&&X<90)&&(Y>90&&Y<100)) || ((X>80&&X<90)&&(Y>90&&Y<140)) || ((X>60&&X<90)&&(Y>130&&Y<140)) || ((X>60&&X<90)&&(Y>110&&Y<120)) ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		else if ((index1==4'd9) && (((X>60&&X<70)&&(Y>90&&Y<120)) || ((X>60&&X<90)&&(Y>90&&Y<100)) || ((X>80&&X<90)&&(Y>90&&Y<140)) || ((X>60&&X<90)&&(Y>110&&Y<120))  ))begin
			colouroutput[11:0] <= 12'b000011111111;
		end
		
		
		
		
		
		else if ( ((X>18 && X<24)&&(Y>169&&Y<181)) || ((X>23&&X<29)&&(Y>179&&Y<191)) || ((X>28&&X<34)&&(Y>189&&Y<201)) || ((X>28&&X<34)&&(Y>149&&Y<201)) || ((X>33&&X<39)&&(Y>179&&Y<191)) || ((X>38&&X<44)&&(Y>169&&Y<181))	)begin// down arrow
			colouroutput[11:0] <= 12'b000011111111;
		end
		//1st character
		else if ((seq2[44:42]==3'b100) &&(((X>20 && X<30)&&(Y>340 && Y<390))||((X>29 && X<50)&&(Y>340 && Y<350))||((X>29 && X<41)&&(Y>365 &&Y<375))||((X>40 && X<50)&&(Y>340 && Y<390)))) begin//"A" at bottom left position
			if (seq2[44:42]==seq1[44:42])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
			end
		else if ((seq2[44:42]==3'b101) && (((X>20 && X<50)&&(Y>340 && Y<350))||((X>20 && X<30)&&(Y>340 && Y<390))||((X>20 && X<50)&&(Y>380 && Y<390))||((X>35 && X<50)&&(Y>360 && Y<370))||((X>40 && X<50)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[44:42]==seq1[44:42])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[44:42]==3'b110) && (((X>20 && X<50)&&(Y>340 && Y<350))||((X>20 && X<30)&&(Y>340 && Y<390))||((X>20 && X<50)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[44:42]==seq1[44:42])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[44:42]==3'b111) && (((X>20&&X<50)&&(Y>340&&Y<350))||((X>30&&X<40)&&(Y>340&&Y<390))))//"T"
			if (seq2[44:42]==seq1[44:42])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[44:42]==3'b010) && (((X>20&&X<50)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;
			
////////////////////////////////////////////////////////////////////////////////			
		else if ((seq2[41:39]==3'b100) &&(((X>60 && X<70)&&(Y>340 && Y<390))||((X>69 && X<90)&&(Y>340 && Y<350))||((X>69 && X<81)&&(Y>365 &&Y<375))||((X>80 && X<90)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[41:39]==seq1[41:39])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[41:39]==3'b101) &&(((X>60 && X<90)&&(Y>340 && Y<350))||((X>60 && X<70)&&(Y>340 && Y<390))||((X>60 && X<90)&&(Y>380 && Y<390))||((X>75 && X<90)&&(Y>360 && Y<370))||((X>80 && X<90)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[41:39]==seq1[41:39])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[41:39]==3'b110) &&(((X>60 && X<90)&&(Y>340 && Y<350))||((X>60 && X<70)&&(Y>340 && Y<390))||((X>60 && X<90)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[41:39]==seq1[41:39])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[41:39]==3'b111) &&(((X>60&&X<90)&&(Y>340&&Y<350))||((X>70&&X<80)&&(Y>340&&Y<390))))//"T"
			if (seq2[41:39]==seq1[41:39])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[41:39]==3'b010) && (((X>60&&X<90)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;
			
			
		else if ((seq2[38:36]==3'b100) &&(((X>100 && X<110)&&(Y>340 && Y<390))||((X>109 && X<130)&&(Y>340 && Y<350))||((X>109 && X<121)&&(Y>365 &&Y<375))||((X>120 && X<130)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[38:36]==seq1[38:36])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[38:36]==3'b101) &&(((X>100 && X<130)&&(Y>340 && Y<350))||((X>100 && X<110)&&(Y>340 && Y<390))||((X>100 && X<130)&&(Y>380 && Y<390))||((X>115 && X<130)&&(Y>360 && Y<370))||((X>120 && X<130)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[38:36]==seq1[38:36])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[38:36]==3'b110) &&(((X>100 && X<130)&&(Y>340 && Y<350))||((X>100 && X<110)&&(Y>340 && Y<390))||((X>100 && X<130)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[38:36]==seq1[38:36])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[38:36]==3'b111) &&(((X>100&&X<130)&&(Y>340&&Y<350))||((X>110&&X<120)&&(Y>340&&Y<390))))//"T"
			if (seq2[38:36]==seq1[38:36])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[38:36]==3'b010) && (((X>100&&X<130)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;
			
			
		else if ((seq2[35:33]==3'b100) &&(((X>140 && X<150)&&(Y>340 && Y<390))||((X>149 && X<170)&&(Y>340 && Y<350))||((X>149 && X<161)&&(Y>365 &&Y<375))||((X>160 && X<170)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[35:33]==seq1[35:33])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[35:33]==3'b101) &&(((X>140 && X<170)&&(Y>340 && Y<350))||((X>140 && X<150)&&(Y>340 && Y<390))||((X>140 && X<170)&&(Y>380 && Y<390))||((X>155 && X<170)&&(Y>360 && Y<370))||((X>160 && X<170)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[35:33]==seq1[35:33])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[35:33]==3'b110) &&(((X>140 && X<170)&&(Y>340 && Y<350))||((X>140 && X<150)&&(Y>340 && Y<390))||((X>140 && X<170)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[35:33]==seq1[35:33])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[35:33]==3'b111) &&(((X>140&&X<170)&&(Y>340&&Y<350))||((X>150&&X<160)&&(Y>340&&Y<390))))//"T"
			if (seq2[35:33]==seq1[35:33])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[35:33]==3'b010) && (((X>140&&X<170)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;
			
			
		else if ((seq2[32:30]==3'b100) &&(((X>180 && X<190)&&(Y>340 && Y<390))||((X>189 && X<210)&&(Y>340 && Y<350))||((X>189 && X<201)&&(Y>365 &&Y<375))||((X>200 && X<210)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[32:30]==seq1[32:30])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[32:30]==3'b101) &&(((X>180 && X<210)&&(Y>340 && Y<350))||((X>180 && X<190)&&(Y>340 && Y<390))||((X>180 && X<210)&&(Y>380 && Y<390))||((X>195 && X<210)&&(Y>360 && Y<370))||((X>200 && X<210)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[32:30]==seq1[32:30])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[32:30]==3'b110) &&(((X>180 && X<210)&&(Y>340 && Y<350))||((X>180 && X<190)&&(Y>340 && Y<390))||((X>180 && X<210)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[32:30]==seq1[32:30])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[32:30]==3'b111) &&(((X>180&&X<210)&&(Y>340&&Y<350))||((X>190&&X<200)&&(Y>340&&Y<390))))//"T"
			if (seq2[32:30]==seq1[32:30])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[32:30]==3'b010) && (((X>180&&X<210)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;	
			
		else if ((seq2[29:27]==3'b100) &&(((X>220 && X<230)&&(Y>340 && Y<390))||((X>229 && X<250)&&(Y>340 && Y<350))||((X>229 && X<241)&&(Y>365 &&Y<375))||((X>240 && X<250)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[29:27]==seq1[29:27])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[29:27]==3'b101) &&(((X>220 && X<250)&&(Y>340 && Y<350))||((X>220 && X<230)&&(Y>340 && Y<390))||((X>220 && X<250)&&(Y>380 && Y<390))||((X>235 && X<250)&&(Y>360 && Y<370))||((X>240 && X<250)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[29:27]==seq1[29:27])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[29:27]==3'b110) &&(((X>220 && X<250)&&(Y>340 && Y<350))||((X>220 && X<230)&&(Y>340 && Y<390))||((X>220 && X<250)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[29:27]==seq1[29:27])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[29:27]==3'b111) &&(((X>220&&X<250)&&(Y>340&&Y<350))||((X>230&&X<240)&&(Y>340&&Y<390))))//"T"
			if (seq2[29:27]==seq1[29:27])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[29:27]==3'b010) && (((X>220&&X<250)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;	
			
			
		else if ((seq2[26:24]==3'b100) &&(((X>260 && X<270)&&(Y>340 && Y<390))||((X>269 && X<290)&&(Y>340 && Y<350))||((X>269 && X<281)&&(Y>365 &&Y<375))||((X>280 && X<290)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[26:24]==seq1[26:24])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[26:24]==3'b101) &&(((X>260 && X<290)&&(Y>340 && Y<350))||((X>260 && X<270)&&(Y>340 && Y<390))||((X>260 && X<290)&&(Y>380 && Y<390))||((X>275 && X<290)&&(Y>360 && Y<370))||((X>280 && X<290)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[26:24]==seq1[26:24])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[26:24]==3'b110) &&(((X>260 && X<290)&&(Y>340 && Y<350))||((X>260 && X<270)&&(Y>340 && Y<390))||((X>260 && X<290)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[26:24]==seq1[26:24])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[26:24]==3'b111) &&(((X>260&&X<290)&&(Y>340&&Y<350))||((X>270&&X<280)&&(Y>340&&Y<390))))//"T"
			if (seq2[26:24]==seq1[26:24])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[26:24]==3'b010) && (((X>260&&X<290)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;	
			
			
		else if ((seq2[23:21]==3'b100) &&(((X>300 && X<310)&&(Y>340 && Y<390))||((X>309 && X<330)&&(Y>340 && Y<350))||((X>309 && X<321)&&(Y>365 &&Y<375))||((X>320 && X<330)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[23:21]==seq1[23:21])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[23:21]==3'b101) &&(((X>300 && X<330)&&(Y>340 && Y<350))||((X>300 && X<310)&&(Y>340 && Y<390))||((X>300 && X<330)&&(Y>380 && Y<390))||((X>315 && X<330)&&(Y>360 && Y<370))||((X>320 && X<330)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[23:21]==seq1[23:21])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[23:21]==3'b110) &&(((X>300 && X<330)&&(Y>340 && Y<350))||((X>300 && X<310)&&(Y>340 && Y<390))||((X>300 && X<330)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[23:21]==seq1[23:21])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[23:21]==3'b111) &&(((X>300&&X<330)&&(Y>340&&Y<350))||((X>310&&X<320)&&(Y>340&&Y<390))))//"T"
			if (seq2[23:21]==seq1[23:21])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[23:21]==3'b010) && (((X>300&&X<330)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;	
			
			
		else if ((seq2[20:18]==3'b100) &&(((X>340 && X<350)&&(Y>340 && Y<390))||((X>349 && X<370)&&(Y>340 && Y<350))||((X>349 && X<361)&&(Y>365 &&Y<375))||((X>360 && X<370)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[20:18]==seq1[20:18])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[20:18]==3'b101) &&(((X>340 && X<370)&&(Y>340 && Y<350))||((X>340 && X<350)&&(Y>340 && Y<390))||((X>340 && X<370)&&(Y>380 && Y<390))||((X>355 && X<370)&&(Y>360 && Y<370))||((X>360 && X<370)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[20:18]==seq1[20:18])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[20:18]==3'b110) &&(((X>340 && X<370)&&(Y>340 && Y<350))||((X>340 && X<350)&&(Y>340 && Y<390))||((X>340 && X<370)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[20:18]==seq1[20:18])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[20:18]==3'b111) &&(((X>340&&X<370)&&(Y>340&&Y<350))||((X>350&&X<360)&&(Y>340&&Y<390))))//"T"
			if (seq2[20:18]==seq1[20:18])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[20:18]==3'b010) && (((X>340&&X<370)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;
			
			
		else if ((seq2[17:15]==3'b100) &&(((X>380 && X<390)&&(Y>340 && Y<390))||((X>389 && X<410)&&(Y>340 && Y<350))||((X>389 && X<401)&&(Y>365 &&Y<375))||((X>400 && X<410)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[17:15]==seq1[17:15])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[17:15]==3'b101) &&(((X>380 && X<410)&&(Y>340 && Y<350))||((X>380 && X<390)&&(Y>340 && Y<390))||((X>380 && X<410)&&(Y>380 && Y<390))||((X>395 && X<410)&&(Y>360 && Y<370))||((X>400 && X<410)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[17:15]==seq1[17:15])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[17:15]==3'b110) &&(((X>380 && X<410)&&(Y>340 && Y<350))||((X>380 && X<390)&&(Y>340 && Y<390))||((X>380 && X<410)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[17:15]==seq1[17:15])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[17:15]==3'b111) &&(((X>380&&X<410)&&(Y>340&&Y<350))||((X>390&&X<400)&&(Y>340&&Y<390))))//"T"
			if (seq2[17:15]==seq1[17:15])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[17:15]==3'b010) && (((X>380&&X<410)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;
			
			
		else if ((seq2[14:12]==3'b100) &&(((X>420 && X<430)&&(Y>340 && Y<390))||((X>429 && X<450)&&(Y>340 && Y<350))||((X>429 && X<441)&&(Y>365 &&Y<375))||((X>440 && X<450)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[14:12]==seq1[14:12])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[14:12]==3'b101) &&(((X>420 && X<450)&&(Y>340 && Y<350))||((X>420 && X<430)&&(Y>340 && Y<390))||((X>420 && X<450)&&(Y>380 && Y<390))||((X>435 && X<450)&&(Y>360 && Y<370))||((X>440 && X<450)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[14:12]==seq1[14:12])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[14:12]==3'b110) &&(((X>420 && X<450)&&(Y>340 && Y<350))||((X>420 && X<430)&&(Y>340 && Y<390))||((X>420 && X<450)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[14:12]==seq1[14:12])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[14:12]==3'b111) &&(((X>420&&X<450)&&(Y>340&&Y<350))||((X>430&&X<440)&&(Y>340&&Y<390))))//"T"
			if (seq2[14:12]==seq1[14:12])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[14:12]==3'b010) && (((X>420&&X<450)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;	
			
			
		else if ((seq2[11:9]==3'b100) &&(((X>460 && X<470)&&(Y>340 && Y<390))||((X>469 && X<490)&&(Y>340 && Y<350))||((X>469 && X<481)&&(Y>365 &&Y<375))||((X>480 && X<490)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[11:9]==seq1[11:9])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[11:9]==3'b101) &&(((X>460 && X<490)&&(Y>340 && Y<350))||((X>460 && X<470)&&(Y>340 && Y<390))||((X>460 && X<490)&&(Y>380 && Y<390))||((X>475 && X<490)&&(Y>360 && Y<370))||((X>480 && X<490)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[11:9]==seq1[11:9])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[11:9]==3'b110) &&(((X>460 && X<490)&&(Y>340 && Y<350))||((X>460 && X<470)&&(Y>340 && Y<390))||((X>460 && X<490)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[11:9]==seq1[11:9])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[11:9]==3'b111) &&(((X>460&&X<490)&&(Y>340&&Y<350))||((X>470&&X<480)&&(Y>340&&Y<390))))//"T"
			if (seq2[11:9]==seq1[11:9])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[11:9]==3'b010) && (((X>460&&X<490)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;		
			
			
		else if ((seq2[8:6]==3'b100) &&(((X>500 && X<510)&&(Y>340 && Y<390))||((X>509 && X<530)&&(Y>340 && Y<350))||((X>509 && X<521)&&(Y>365 &&Y<375))||((X>520 && X<530)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[8:6]==seq1[8:6])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[8:6]==3'b101) &&(((X>500 && X<530)&&(Y>340 && Y<350))||((X>500 && X<510)&&(Y>340 && Y<390))||((X>500 && X<530)&&(Y>380 && Y<390))||((X>515 && X<530)&&(Y>360 && Y<370))||((X>520 && X<530)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[8:6]==seq1[8:6])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[8:6]==3'b110) &&(((X>500 && X<530)&&(Y>340 && Y<350))||((X>500 && X<510)&&(Y>340 && Y<390))||((X>500 && X<530)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[8:6]==seq1[8:6])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[8:6]==3'b111) &&(((X>500&&X<530)&&(Y>340&&Y<350))||((X>510&&X<520)&&(Y>340&&Y<390))))//"T"
			if (seq2[8:6]==seq1[8:6])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[8:6]==3'b010) && (((X>500&&X<530)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;		


		else if ((seq2[5:3]==3'b100) &&(((X>540 && X<550)&&(Y>340 && Y<390))||((X>549 && X<570)&&(Y>340 && Y<350))||((X>549 && X<561)&&(Y>365 &&Y<375))||((X>560 && X<570)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[5:3]==seq1[5:3])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[5:3]==3'b101) &&(((X>540 && X<570)&&(Y>340 && Y<350))||((X>540 && X<550)&&(Y>340 && Y<390))||((X>540 && X<570)&&(Y>380 && Y<390))||((X>555 && X<570)&&(Y>360 && Y<370))||((X>560 && X<570)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[5:3]==seq1[5:3])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[5:3]==3'b110) &&(((X>540 && X<570)&&(Y>340 && Y<350))||((X>540 && X<550)&&(Y>340 && Y<390))||((X>540 && X<570)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[5:3]==seq1[5:3])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[5:3]==3'b111) &&(((X>540&&X<570)&&(Y>340&&Y<350))||((X>550&&X<560)&&(Y>340&&Y<390))))//"T"
			if (seq2[5:3]==seq1[5:3])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[5:3]==3'b010) && (((X>540&&X<570)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;				
	
	
		else if ((seq2[2:0]==3'b100) &&(((X>580 && X<590)&&(Y>340 && Y<390))||((X>589 && X<610)&&(Y>340 && Y<350))||((X>589 && X<601)&&(Y>365 &&Y<375))||((X>600 && X<610)&&(Y>340 && Y<390)))) //"A" at bottom left position
			if (seq2[2:0]==seq1[2:0])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[2:0]==3'b101) &&(((X>580 && X<610)&&(Y>340 && Y<350))||((X>580 && X<590)&&(Y>340 && Y<390))||((X>580 && X<610)&&(Y>380 && Y<390))||((X>595 && X<610)&&(Y>360 && Y<370))||((X>600 && X<610)&&(Y>360 && Y<390))))//"G" beside A 
			if (seq2[2:0]==seq1[2:0])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[2:0]==3'b110) &&(((X>580 && X<610)&&(Y>340 && Y<350))||((X>580 && X<590)&&(Y>340 && Y<390))||((X>580 && X<610)&&(Y>380 && Y<390))))//"G" beside A 
			if (seq2[2:0]==seq1[2:0])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[2:0]==3'b111) &&(((X>580&&X<610)&&(Y>340&&Y<350))||((X>590&&X<600)&&(Y>340&&Y<390))))//"T"
			if (seq2[2:0]==seq1[2:0])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq2[2:0]==3'b010) && (((X>580&&X<610)&&(Y>360&&Y<370))))//"-"
			colouroutput[11:0]<= 12'b111100000000;		
			//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
			//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
			//seq1
			
		else if ((seq1[44:42]==3'b100) &&(((X>20 && X<30)&&(Y>210 && Y<260))||((X>20 && X<50)&&(Y>210 && Y<220))||((X>40 && X<50)&&(Y>210 && Y<260))||((X>29 && X<41)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[44:42]==seq1[44:42])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[44:42]==3'b101) &&(((X>20 && X<50)&&(Y>210 && Y<220))||((X>20 && X<30)&&(Y>210 && Y<260))||((X>20 && X<50)&&(Y>250 && Y<260))||((X>40 && X<50)&&(Y>230 && Y<260))||((X>45 && X<50)&&(Y>230 && Y<240))))//"G" 
			if (seq2[44:42]==seq1[44:42])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[44:42]==3'b110) &&(((X>20 && X<50)&&(Y>210 && Y<220))||((X>20 && X<30)&&(Y>210 && Y<260))||((X>20 && X<50)&&(Y>250 && Y<260))))//"C" 
			if (seq2[44:42]==seq1[44:42])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[44:42]==3'b111) &&(((X>20&&X<50)&&(Y>210&&Y<220))||((X>30&&X<40)&&(Y>210&&Y<260))))//"T"
			if (seq2[44:42]==seq1[44:42])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[44:42]==3'b010) && ((X>20&&X<50)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;
		
		///////////////////////////////////////

		else if ((seq1[41:39]==3'b100) &&(((X>60 && X<70)&&(Y>210 && Y<260))||((X>60 && X<90)&&(Y>210 && Y<220))||((X>80 && X<90)&&(Y>210 && Y<260))||((X>69 && X<81)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[41:39]==seq1[41:39])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[41:39]==3'b101) &&(((X>60 && X<90)&&(Y>210 && Y<220))||((X>60 && X<70)&&(Y>210 && Y<260))||((X>60 && X<90)&&(Y>250 && Y<260))||((X>80 && X<90)&&(Y>230 && Y<260))||((X>85 && X<90)&&(Y>230 && Y<240))))//"G" 
			if (seq2[41:39]==seq1[41:39])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[41:39]==3'b110) &&(((X>60 && X<90)&&(Y>210 && Y<220))||((X>60 && X<70)&&(Y>210 && Y<260))||((X>60 && X<90)&&(Y>250 && Y<260))))//"C" 
			if (seq2[41:39]==seq1[41:39])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[41:39]==3'b111) &&(((X>60&&X<90)&&(Y>210&&Y<220))||((X>70&&X<80)&&(Y>210&&Y<260))))//"T"
			if (seq2[41:39]==seq1[41:39])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[41:39]==3'b010) && ((X>60&&X<90)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;
		
		////////////////////////////////////////////
		
		else if ((seq1[38:36]==3'b100) &&(((X>100 && X<110)&&(Y>210 && Y<260))||((X>100 && X<130)&&(Y>210 && Y<220))||((X>120 && X<130)&&(Y>210 && Y<260))||((X>109 && X<121)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[38:36]==seq1[38:36])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[38:36]==3'b101) &&(((X>100 && X<130)&&(Y>210 && Y<220))||((X>100 && X<110)&&(Y>210 && Y<260))||((X>100 && X<130)&&(Y>250 && Y<260))||((X>120 && X<130)&&(Y>230 && Y<260))||((X>125 && X<130)&&(Y>230 && Y<240))))//"G" 
			if (seq2[38:36]==seq1[38:36])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[38:36]==3'b110) &&(((X>100 && X<130)&&(Y>210 && Y<220))||((X>100 && X<110)&&(Y>210 && Y<260))||((X>100 && X<130)&&(Y>250 && Y<260))))//"C" 
			if (seq2[38:36]==seq1[38:36])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[38:36]==3'b111) &&(((X>100&&X<130)&&(Y>210&&Y<220))||((X>110&&X<120)&&(Y>210&&Y<260))))//"T"
			if (seq2[38:36]==seq1[38:36])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[38:36]==3'b010) && ((X>100&&X<130)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;
		
		////////////////////////////////////////////
			
		else if ((seq1[35:33]==3'b100) &&(((X>140 && X<150)&&(Y>210 && Y<260))||((X>140 && X<170)&&(Y>210 && Y<220))||((X>160 && X<170)&&(Y>210 && Y<260))||((X>149 && X<161)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[35:33]==seq1[35:33])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[35:33]==3'b101) &&(((X>140 && X<170)&&(Y>210 && Y<220))||((X>140 && X<150)&&(Y>210 && Y<260))||((X>140 && X<170)&&(Y>250 && Y<260))||((X>160 && X<170)&&(Y>230 && Y<260))||((X>165 && X<170)&&(Y>230 && Y<240))))//"G" 
			if (seq2[35:33]==seq1[35:33])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[35:33]==3'b110) &&(((X>140 && X<170)&&(Y>210 && Y<220))||((X>140 && X<150)&&(Y>210 && Y<260))||((X>140 && X<170)&&(Y>250 && Y<260))))//"C" 
			if (seq2[35:33]==seq1[35:33])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[35:33]==3'b111) &&(((X>140&&X<170)&&(Y>210&&Y<220))||((X>150&&X<160)&&(Y>210&&Y<260))))//"T"
			if (seq2[35:33]==seq1[35:33])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[35:33]==3'b010) && ((X>140&&X<170)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;
		
		////////////////////////////////////////////	
		
		else if ((seq1[32:30]==3'b100) &&(((X>180 && X<190)&&(Y>210 && Y<260))||((X>180 && X<210)&&(Y>210 && Y<220))||((X>200 && X<210)&&(Y>210 && Y<260))||((X>189 && X<201)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[32:30]==seq1[32:30])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[32:30]==3'b101) &&(((X>180 && X<210)&&(Y>210 && Y<220))||((X>180 && X<190)&&(Y>210 && Y<260))||((X>180 && X<210)&&(Y>250 && Y<260))||((X>200 && X<210)&&(Y>230 && Y<260))||((X>205 && X<210)&&(Y>230 && Y<240))))//"G" 
			if (seq2[32:30]==seq1[32:30])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[32:30]==3'b110) &&(((X>180 && X<210)&&(Y>210 && Y<220))||((X>180 && X<190)&&(Y>210 && Y<260))||((X>180 && X<210)&&(Y>250 && Y<260))))//"C" 
			if (seq2[32:30]==seq1[32:30])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[32:30]==3'b111) &&(((X>180&&X<210)&&(Y>210&&Y<220))||((X>190&&X<200)&&(Y>210&&Y<260))))//"T"
			if (seq2[32:30]==seq1[32:30])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[32:30]==3'b010) && ((X>180&&X<210)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;
		
		////////////////////////////////////////////
			
		else if ((seq1[29:27]==3'b100) &&(((X>220 && X<230)&&(Y>210 && Y<260))||((X>220 && X<250)&&(Y>210 && Y<220))||((X>240 && X<250)&&(Y>210 && Y<260))||((X>229 && X<241)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[29:27]==seq1[29:27])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[29:27]==3'b101) &&(((X>220 && X<250)&&(Y>210 && Y<220))||((X>220 && X<230)&&(Y>210 && Y<260))||((X>220 && X<250)&&(Y>250 && Y<260))||((X>240 && X<250)&&(Y>230 && Y<260))||((X>245 && X<250)&&(Y>230 && Y<240))))//"G" 
			if (seq2[29:27]==seq1[29:27])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[29:27]==3'b110) &&(((X>220 && X<250)&&(Y>210 && Y<220))||((X>220 && X<230)&&(Y>210 && Y<260))||((X>220 && X<250)&&(Y>250 && Y<260))))//"C" 
			if (seq2[29:27]==seq1[29:27])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[29:27]==3'b111) &&(((X>220&&X<250)&&(Y>210&&Y<220))||((X>230&&X<240)&&(Y>210&&Y<260))))//"T"
			if (seq2[29:27]==seq1[29:27])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[29:27]==3'b010) && ((X>220&&X<250)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;
		
		////////////////////////////////////////////

		else if ((seq1[26:24]==3'b100) &&(((X>260 && X<270)&&(Y>210 && Y<260))||((X>260 && X<290)&&(Y>210 && Y<220))||((X>280 && X<290)&&(Y>210 && Y<260))||((X>269 && X<281)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[26:24]==seq1[26:24])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[26:24]==3'b101) &&(((X>260 && X<290)&&(Y>210 && Y<220))||((X>260 && X<270)&&(Y>210 && Y<260))||((X>260 && X<290)&&(Y>250 && Y<260))||((X>280 && X<290)&&(Y>230 && Y<260))||((X>285 && X<290)&&(Y>230 && Y<240))))//"G" 
			if (seq2[26:24]==seq1[26:24])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[26:24]==3'b110) &&(((X>260 && X<290)&&(Y>210 && Y<220))||((X>260 && X<270)&&(Y>210 && Y<260))||((X>260 && X<290)&&(Y>250 && Y<260))))//"C" 
			if (seq2[26:24]==seq1[26:24])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[26:24]==3'b111) &&(((X>260&&X<290)&&(Y>210&&Y<220))||((X>270&&X<280)&&(Y>210&&Y<260))))//"T"
			if (seq2[26:24]==seq1[26:24])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[26:24]==3'b010) && ((X>260&&X<290)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;
		
		////////////////////////////////////////////
		
		else if ((seq1[23:21]==3'b100) &&(((X>300 && X<310)&&(Y>210 && Y<260))||((X>300 && X<330)&&(Y>210 && Y<220))||((X>320 && X<330)&&(Y>210 && Y<260))||((X>309 && X<321)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[23:21]==seq1[23:21])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[23:21]==3'b101) &&(((X>300 && X<330)&&(Y>210 && Y<220))||((X>300 && X<310)&&(Y>210 && Y<260))||((X>300 && X<330)&&(Y>250 && Y<260))||((X>320 && X<330)&&(Y>230 && Y<260))||((X>325 && X<330)&&(Y>230 && Y<240))))//"G" 
			if (seq2[23:21]==seq1[23:21])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[23:21]==3'b110) &&(((X>300 && X<330)&&(Y>210 && Y<220))||((X>300 && X<310)&&(Y>210 && Y<260))||((X>300 && X<330)&&(Y>250 && Y<260))))//"C" 
			if (seq2[23:21]==seq1[23:21])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[23:21]==3'b111) &&(((X>300&&X<330)&&(Y>210&&Y<220))||((X>310&&X<320)&&(Y>210&&Y<260))))//"T"
			if (seq2[23:21]==seq1[23:21])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[23:21]==3'b010) && ((X>300&&X<330)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;
		
		else if ((seq1[20:18]==3'b100) &&(((X>340 && X<350)&&(Y>210 && Y<260))||((X>340 && X<370)&&(Y>210 && Y<220))||((X>360 && X<370)&&(Y>210 && Y<260))||((X>349 && X<361)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[20:18]==seq1[20:18])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[20:18]==3'b101) &&(((X>340 && X<370)&&(Y>210 && Y<220))||((X>340 && X<350)&&(Y>210 && Y<260))||((X>340 && X<370)&&(Y>250 && Y<260))||((X>360 && X<370)&&(Y>230 && Y<260))||((X>365 && X<370)&&(Y>230 && Y<240))))//"G" 
			if (seq2[20:18]==seq1[20:18])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[20:18]==3'b110) &&(((X>340 && X<370)&&(Y>210 && Y<220))||((X>340 && X<350)&&(Y>210 && Y<260))||((X>340 && X<370)&&(Y>250 && Y<260))))//"C" 
			if (seq2[20:18]==seq1[20:18])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[20:18]==3'b111) &&(((X>340&&X<370)&&(Y>210&&Y<220))||((X>350&&X<360)&&(Y>210&&Y<260))))//"T"
			if (seq2[20:18]==seq1[20:18])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[20:18]==3'b010) && ((X>340&&X<370)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;
			
		else if ((seq1[17:15]==3'b100) &&(((X>380 && X<390)&&(Y>210 && Y<260))||((X>380 && X<410)&&(Y>210 && Y<220))||((X>400 && X<410)&&(Y>210 && Y<260))||((X>389 && X<401)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[17:15]==seq1[17:15])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[17:15]==3'b101) &&(((X>380 && X<410)&&(Y>210 && Y<220))||((X>380 && X<390)&&(Y>210 && Y<260))||((X>380 && X<410)&&(Y>250 && Y<260))||((X>400 && X<410)&&(Y>230 && Y<260))||((X>405 && X<410)&&(Y>230 && Y<240))))//"G" 
			if (seq2[17:15]==seq1[17:15])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[17:15]==3'b110) &&(((X>380 && X<410)&&(Y>210 && Y<220))||((X>380 && X<390)&&(Y>210 && Y<260))||((X>380 && X<410)&&(Y>250 && Y<260))))//"C" 
			if (seq2[17:15]==seq1[17:15])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[17:15]==3'b111) &&(((X>380&&X<410)&&(Y>210&&Y<220))||((X>390&&X<400)&&(Y>210&&Y<260))))//"T"
			if (seq2[17:15]==seq1[17:15])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[17:15]==3'b010) && ((X>380&&X<410)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;		
	
		else if ((seq1[14:12]==3'b100) &&(((X>420 && X<430)&&(Y>210 && Y<260))||((X>420 && X<450)&&(Y>210 && Y<220))||((X>440 && X<450)&&(Y>210 && Y<260))||((X>429 && X<441)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[14:12]==seq1[14:12])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[14:12]==3'b101) &&(((X>420 && X<450)&&(Y>210 && Y<220))||((X>420 && X<430)&&(Y>210 && Y<260))||((X>420 && X<450)&&(Y>250 && Y<260))||((X>440 && X<450)&&(Y>230 && Y<260))||((X>445 && X<450)&&(Y>230 && Y<240))))//"G" 
			if (seq2[14:12]==seq1[14:12])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[14:12]==3'b110) &&(((X>420 && X<450)&&(Y>210 && Y<220))||((X>420 && X<430)&&(Y>210 && Y<260))||((X>420 && X<450)&&(Y>250 && Y<260))))//"C" 
			if (seq2[14:12]==seq1[14:12])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[14:12]==3'b111) &&(((X>420&&X<450)&&(Y>210&&Y<220))||((X>430&&X<440)&&(Y>210&&Y<260))))//"T"
			if (seq2[14:12]==seq1[14:12])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[14:12]==3'b010) && ((X>420&&X<450)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;	
		
		else if ((seq1[11:9]==3'b100) &&(((X>460 && X<470)&&(Y>210 && Y<260))||((X>460 && X<490)&&(Y>210 && Y<220))||((X>480 && X<490)&&(Y>210 && Y<260))||((X>469 && X<481)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[11:9]==seq1[11:9])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[11:9]==3'b101) &&(((X>460 && X<490)&&(Y>210 && Y<220))||((X>460 && X<470)&&(Y>210 && Y<260))||((X>460 && X<490)&&(Y>250 && Y<260))||((X>480 && X<490)&&(Y>230 && Y<260))||((X>485 && X<490)&&(Y>230 && Y<240))))//"G" 
			if (seq2[11:9]==seq1[11:9])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[11:9]==3'b110) &&(((X>460 && X<490)&&(Y>210 && Y<220))||((X>460 && X<470)&&(Y>210 && Y<260))||((X>460 && X<490)&&(Y>250 && Y<260))))//"C" 
			if (seq2[11:9]==seq1[11:9])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[11:9]==3'b111) &&(((X>460&&X<490)&&(Y>210&&Y<220))||((X>470&&X<480)&&(Y>210&&Y<260))))//"T"
			if (seq2[11:9]==seq1[11:9])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[11:9]==3'b010) && ((X>460&&X<490)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;			
	
		else if ((seq1[8:6]==3'b100) &&(((X>500 && X<510)&&(Y>210 && Y<260))||((X>500 && X<530)&&(Y>210 && Y<220))||((X>520 && X<530)&&(Y>210 && Y<260))||((X>509 && X<521)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[8:6]==seq1[8:6])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[8:6]==3'b101) &&(((X>500 && X<530)&&(Y>210 && Y<220))||((X>500 && X<510)&&(Y>210 && Y<260))||((X>500 && X<530)&&(Y>250 && Y<260))||((X>520 && X<530)&&(Y>230 && Y<260))||((X>525 && X<530)&&(Y>230 && Y<240))))//"G" 
			if (seq2[8:6]==seq1[8:6])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[8:6]==3'b110) &&(((X>500 && X<530)&&(Y>210 && Y<220))||((X>500 && X<510)&&(Y>210 && Y<260))||((X>500 && X<530)&&(Y>250 && Y<260))))//"C" 
			if (seq2[8:6]==seq1[8:6])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[8:6]==3'b111) &&(((X>500&&X<530)&&(Y>210&&Y<220))||((X>510&&X<520)&&(Y>210&&Y<260))))//"T"
			if (seq2[8:6]==seq1[8:6])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[8:6]==3'b010) && ((X>500&&X<530)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;	

		else if ((seq1[5:3]==3'b100) &&(((X>540 && X<550)&&(Y>210 && Y<260))||((X>540 && X<570)&&(Y>210 && Y<220))||((X>560 && X<570)&&(Y>210 && Y<260))||((X>549 && X<561)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[5:3]==seq1[5:3])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[5:3]==3'b101) &&(((X>540 && X<570)&&(Y>210 && Y<220))||((X>540 && X<550)&&(Y>210 && Y<260))||((X>540 && X<570)&&(Y>250 && Y<260))||((X>560 && X<570)&&(Y>230 && Y<260))||((X>565 && X<570)&&(Y>230 && Y<240))))//"G" 
			if (seq2[5:3]==seq1[5:3])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[5:3]==3'b110) &&(((X>540 && X<570)&&(Y>210 && Y<220))||((X>540 && X<550)&&(Y>210 && Y<260))||((X>540 && X<570)&&(Y>250 && Y<260))))//"C" 
			if (seq2[5:3]==seq1[5:3])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[5:3]==3'b111) &&(((X>540&&X<570)&&(Y>210&&Y<220))||((X>550&&X<560)&&(Y>210&&Y<260))))//"T"
			if (seq2[5:3]==seq1[5:3])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[5:3]==3'b010) && ((X>540&&X<570)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;

		else if ((seq1[2:0]==3'b100) &&(((X>580 && X<590)&&(Y>210 && Y<260))||((X>580 && X<610)&&(Y>210 && Y<220))||((X>600 && X<610)&&(Y>210 && Y<260))||((X>589 && X<601)&&(Y>235 && Y<245)))) //"A" 
			if (seq2[2:0]==seq1[2:0])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[2:0]==3'b101) &&(((X>580 && X<610)&&(Y>210 && Y<220))||((X>580 && X<590)&&(Y>210 && Y<260))||((X>580 && X<610)&&(Y>250 && Y<260))||((X>600 && X<610)&&(Y>230 && Y<260))||((X>605 && X<610)&&(Y>230 && Y<240))))//"G" 
			if (seq2[2:0]==seq1[2:0])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[2:0]==3'b110) &&(((X>580 && X<610)&&(Y>210 && Y<220))||((X>580 && X<590)&&(Y>210 && Y<260))||((X>580 && X<610)&&(Y>250 && Y<260))))//"C" 
			if (seq2[2:0]==seq1[2:0])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[2:0]==3'b111) &&(((X>580&&X<610)&&(Y>210&&Y<220))||((X>590&&X<600)&&(Y>210&&Y<260))))//"T"
			if (seq2[2:0]==seq1[2:0])
				colouroutput[11:0]<= 12'b000011110000;
			else
				colouroutput[11:0]<= 12'b111100000000;
		else if ((seq1[2:0]==3'b010) && ((X>580&&X<610)&&(Y>230&&Y<240)))//"___"
			colouroutput[11:0]<= 12'b111100000000;	
	
		else 
			colouroutput[11:0]<= 12'b011101110111;
			//colouroutput[11:0]<= 12'b000000000000;
	end
end	
assign VGA_R = colouroutput[11:8];
assign VGA_G = colouroutput[7:4];
assign VGA_B = colouroutput[3:0];

endmodule